module adder;

endmodule

// adder