module data_memory;

endmodule

// data_memory