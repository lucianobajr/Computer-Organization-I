module alu;

endmodule

// alu