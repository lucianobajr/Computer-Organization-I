module sign_extended;

endmodule

// sign_extended