// ADD, SUB, AND, OR, LD, SD, BEQ

module main;

endmodule

// Main