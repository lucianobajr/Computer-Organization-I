module intruction_memory;

endmodule

// intruction_memory