module imm_gen;

endmodule

// imm_gen