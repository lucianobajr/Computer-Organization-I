module mux;

endmodule

// mux