module pc;

endmodule

// pc