module reg_file;

endmodule

// reg_file