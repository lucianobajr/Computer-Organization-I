module controle;

endmodule

// control